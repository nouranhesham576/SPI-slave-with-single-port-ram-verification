interface SPI_Wrapper_interface (input bit clk);
logic rst_n;
logic MOSI;
logic MISO;
logic SS_n;
logic MISO_golden;



endinterface