package SPI_shared_pkg;
    bit[5:0] count;
    logic [10:0] arr_of_data;
    bit is_read;
    bit have_address_to_read;
    int limit;
endpackage